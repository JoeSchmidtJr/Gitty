module test;
    initial begin
        $display("HEY WHAT.");
        $finish;
    end
endmodule